`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08/06/2025 04:22:54 PM
// Design Name: 
// Module Name: Swap_FSM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Swap_FSM(
input clk , reset_n,swap,
output we ,
input [1:0] sel);

reg [1:0] state_reg , state_next;
parameter s0=0 , s1=1 , s2=2 , s3=3 ;
//current state logic
always@(posedge clk , negedge reset_n)
begin
    if(~reset_n)
    state_reg <= 'b0;
    else
    state_reg <= state_next;
end
//Next state logic
always@(*)
begin
    case(state_reg)
     s0: if(~swap)
            state_next = s0 ;
         else
            state_next = s1 ;
     s1: state_next = s2 ;
     s2: state_next = s3 ;
     s3: state_next = s0 ;
default: state_next = s0 ;
    endcase
end

// Output logic
assign sel =  state_reg ;
assign we  = ( state_reg != s0) ;

endmodule
